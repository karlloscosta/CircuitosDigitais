module comparador();
    logic aeqb;
    logic altb;
    logic agtb;

comparador comparador( 
    .aeqb(aeqb),
    .altb(altb),
    .agtb(agtb)
);


endmodule
